//include "core_defines.vh"

module dcache(
  input clock, reset
);

endmodule