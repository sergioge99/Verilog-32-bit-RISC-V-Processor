//include "core_defines.vh"

module mul(
  input clock, reset
);

endmodule