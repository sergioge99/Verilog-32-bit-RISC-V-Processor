//include "core_defines.vh"

module C_top(
  input clock, reset
);

endmodule
