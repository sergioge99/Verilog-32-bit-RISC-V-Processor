//include "core_defines.vh"

module itlb(
  input clock, reset
);

endmodule
