//include "core_defines.vh"

module alu(
  input clock, reset
);

endmodule