//include "core_defines.vh"

module regfile(
  input clock, reset
);

endmodule