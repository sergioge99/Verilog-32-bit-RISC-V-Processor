//include "core_defines.vh"

module dtlb(
  input clock, reset
);

endmodule