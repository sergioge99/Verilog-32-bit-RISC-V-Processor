//include "core_defines.vh"

module A_top(
  input clock, reset
);

endmodule
