//include "core_defines.vh"

module decoder(
  input clock, reset
);

endmodule