//include "core_defines.vh"

module ROB(
  input clock, reset
);

endmodule
