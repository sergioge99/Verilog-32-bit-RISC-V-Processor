//include "core_defines.vh"

module W_top(
  input clock, reset
);

endmodule
