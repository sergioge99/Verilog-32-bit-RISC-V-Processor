//include "core_defines.vh"

module icache(
  input clock, reset,
  input [31:0] addr, 
  output [31:0] instr
);

reg [31:0] icache[31:0];//32 instrucciones de 32 bits de momento

initial begin
  //Aqui se leerá de un fichero las instr
  //pero de momento...
  icache[0] <= 32'h3e800093;
  icache[1] <= 32'h7d008113;
  icache[2] <= 32'hc1810193;
  icache[3] <= 32'h83018213;
  icache[4] <= 32'h3e820293;
  icache[5] <= 32'b00000000000000000000000000000000;
  icache[6] <= 32'b00000000000000000000000000000000;
  icache[7] <= 32'b00000000000000000000000000000000;
  icache[8] <= 32'b00000000000000000000000000000000;
  icache[9] <= 32'b00000000000000000000000000000000;
  icache[10] <= 32'b00000000000000000000000000000000;
  icache[11] <= 32'b00000000000000000000000000000000;
  icache[12] <= 32'b00000000000000000000000000000000;
  icache[13] <= 32'b00000000000000000000000000000000;
  icache[14] <= 32'b00000000000000000000000000000000;
  icache[15] <= 32'b00000000000000000000000000000000;
  icache[16] <= 32'b00000000000000000000000000000000;
  icache[17] <= 32'b00000000000000000000000000000000;
  icache[18] <= 32'b00000000000000000000000000000000;
  icache[19] <= 32'b00000000000000000000000000000000;
  icache[20] <= 32'b00000000000000000000000000000000;
  icache[21] <= 32'b00000000000000000000000000000000;
end

assign instr = icache[addr/4];


endmodule